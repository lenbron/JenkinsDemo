module demo;
	
	initial begin
		$display("Hello world111!!!!");
	end
endmodule
