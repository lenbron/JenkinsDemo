module demo;
	
	initial begin
		$display("Hello world1!!!!");
	end
endmodule
