module demo;
	
	initial begin
		$display("Hello world!!!!");
	end
endmodule
