module demo;
	
	initial begin
		$display("Hello world1111111!!!!");
	end
endmodule
